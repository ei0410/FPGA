`timescale 1ns / 1ps

module led(s1, q);
	input  wire s1;
	output wire q;
	
	assign q = s1;
endmodule
